library verilog;
use verilog.vl_types.all;
entity somador8_vlg_vec_tst is
end somador8_vlg_vec_tst;
